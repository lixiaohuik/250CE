module CE(input clk, input reset,
    input [39:0] io_signalIn_real,
    input [39:0] io_signalIn_imag,
    output[39:0] io_signalOut_real,
    output[39:0] io_signalOut_imag
);

  wire[39:0] T0;
  wire[39:0] T1;
  wire[39:0] T236;
  wire[40:0] T2;
  wire[40:0] T3;
  wire[40:0] T237;
  wire[64:0] T4;
  wire[64:0] T5;
  wire[64:0] T238;
  wire[40:0] T6;
  wire[40:0] T7;
  wire[72:0] T8;
  wire[72:0] T239;
  wire[79:0] T9;
  wire[39:0] T10;
  wire[39:0] T11;
  wire[39:0] T12;
  wire[33:0] T13;
  wire[33:0] T14;
  reg [33:0] stored_Weight_i_0;
  wire[33:0] T240;
  wire[33:0] T15;
  wire[33:0] T16;
  wire[33:0] T241;
  wire[46:0] T17;
  wire[46:0] T18;
  wire[46:0] T242;
  wire[64:0] T19;
  wire[64:0] T20;
  wire[64:0] T243;
  wire[46:0] T21;
  wire[46:0] T22;
  wire[78:0] T23;
  wire[78:0] T244;
  wire[79:0] T24;
  wire[79:0] T25;
  wire[79:0] T26;
  wire[79:0] T27;
  wire[79:0] T28;
  wire[78:0] T29;
  wire[78:0] T30;
  wire[78:0] T245;
  wire[81:0] T31;
  wire[40:0] T32;
  wire[40:0] T33;
  wire[39:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire[40:0] T38;
  wire[40:0] T39;
  wire[40:0] T40;
  wire[40:0] T41;
  wire[40:0] T42;
  wire[40:0] T43;
  wire[40:0] T44;
  wire[40:0] T45;
  wire[39:0] T46;
  wire T47;
  wire T48;
  wire T49;
  wire[40:0] T50;
  wire[40:0] T51;
  wire[39:0] T52;
  wire[39:0] T53;
  wire[33:0] T54;
  wire[5:0] T55;
  wire[3:0] T56;
  wire[1:0] T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire[79:0] T65;
  wire[78:0] T66;
  wire[78:0] T67;
  wire[65:0] T68;
  wire[65:0] T69;
  wire[12:0] T70;
  wire[11:0] T71;
  wire[7:0] T72;
  wire[3:0] T73;
  wire[1:0] T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire[17:0] T246;
  wire T247;
  wire T81;
  wire T82;
  wire[1:0] T83;
  reg [33:0] stored_Weight_i_1;
  wire[33:0] T248;
  wire[33:0] T93;
  wire T94;
  wire T95;
  wire T84;
  wire T249;
  reg [31:0] PTCount;
  wire[31:0] T250;
  wire[31:0] T85;
  wire[31:0] T86;
  wire T87;
  wire T88;
  reg [31:0] sigCount;
  wire[31:0] T251;
  wire[31:0] T89;
  wire[31:0] T90;
  wire[31:0] T91;
  wire[31:0] T92;
  wire[5:0] T96;
  wire[3:0] T97;
  wire[1:0] T98;
  wire T99;
  wire T100;
  wire T101;
  wire[23:0] T252;
  wire T253;
  wire[39:0] T102;
  wire[39:0] T254;
  wire[40:0] T103;
  wire[40:0] T104;
  wire[40:0] T255;
  wire[64:0] T105;
  wire[64:0] T106;
  wire[64:0] T256;
  wire[40:0] T107;
  wire[40:0] T108;
  wire[72:0] T109;
  wire[72:0] T257;
  wire[79:0] T110;
  wire[39:0] T111;
  wire[39:0] T112;
  wire[39:0] T113;
  wire[33:0] T114;
  wire[5:0] T115;
  wire[3:0] T116;
  wire[1:0] T117;
  wire T118;
  wire T119;
  wire T120;
  wire[23:0] T258;
  wire T259;
  wire T121;
  wire[1:0] T122;
  wire[39:0] T123;
  wire[39:0] T124;
  wire[39:0] T260;
  wire[40:0] T125;
  wire[40:0] T126;
  wire[40:0] T261;
  wire[64:0] T127;
  wire[64:0] T128;
  wire[64:0] T262;
  wire[40:0] T129;
  wire[40:0] T130;
  wire[72:0] T131;
  wire[72:0] T263;
  wire[79:0] T132;
  wire[39:0] T133;
  wire[39:0] T134;
  wire[39:0] T135;
  wire[33:0] T136;
  wire[33:0] T137;
  reg [33:0] stored_Weight_r_0;
  wire[33:0] T264;
  wire[33:0] T138;
  wire[33:0] T139;
  wire[33:0] T265;
  wire[46:0] T140;
  wire[46:0] T141;
  wire[46:0] T266;
  wire[64:0] T142;
  wire[64:0] T143;
  wire[64:0] T267;
  wire[46:0] T144;
  wire[46:0] T145;
  wire[78:0] T146;
  wire[78:0] T268;
  wire[79:0] T147;
  wire[79:0] T148;
  wire[79:0] T149;
  wire[79:0] T150;
  wire[79:0] T151;
  wire[78:0] T152;
  wire[78:0] T153;
  wire[78:0] T269;
  wire[81:0] T154;
  wire[40:0] T155;
  wire[40:0] T156;
  wire[39:0] T157;
  wire T158;
  wire T159;
  wire T160;
  wire[40:0] T161;
  wire[40:0] T162;
  wire[40:0] T163;
  wire[40:0] T164;
  wire[40:0] T165;
  wire[40:0] T166;
  wire[40:0] T167;
  wire[40:0] T168;
  wire[39:0] T169;
  wire T170;
  wire T171;
  wire T172;
  wire[40:0] T173;
  wire[40:0] T174;
  wire[39:0] T175;
  wire[39:0] T176;
  wire[33:0] T177;
  wire[5:0] T178;
  wire[3:0] T179;
  wire[1:0] T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire[79:0] T188;
  wire[78:0] T189;
  wire[78:0] T190;
  wire[65:0] T191;
  wire[65:0] T192;
  wire[12:0] T193;
  wire[11:0] T194;
  wire[7:0] T195;
  wire[3:0] T196;
  wire[1:0] T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire[17:0] T270;
  wire T271;
  wire T204;
  wire T205;
  wire[1:0] T206;
  reg [33:0] stored_Weight_r_1;
  wire[33:0] T272;
  wire[33:0] T208;
  wire T209;
  wire T210;
  wire T207;
  wire T273;
  wire[5:0] T211;
  wire[3:0] T212;
  wire[1:0] T213;
  wire T214;
  wire T215;
  wire T216;
  wire[23:0] T274;
  wire T275;
  wire[39:0] T217;
  wire[39:0] T276;
  wire[40:0] T218;
  wire[40:0] T219;
  wire[40:0] T277;
  wire[64:0] T220;
  wire[64:0] T221;
  wire[64:0] T278;
  wire[40:0] T222;
  wire[40:0] T223;
  wire[72:0] T224;
  wire[72:0] T279;
  wire[79:0] T225;
  wire[39:0] T226;
  wire[39:0] T227;
  wire[39:0] T228;
  wire[33:0] T229;
  wire[5:0] T230;
  wire[3:0] T231;
  wire[1:0] T232;
  wire T233;
  wire T234;
  wire T235;
  wire[23:0] T280;
  wire T281;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    stored_Weight_i_0 = {2{$random}};
    stored_Weight_i_1 = {2{$random}};
    PTCount = {1{$random}};
    sigCount = {1{$random}};
    stored_Weight_r_0 = {2{$random}};
    stored_Weight_r_1 = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_signalOut_imag = T0;
  assign T0 = T121 ? T102 : T1;
  assign T1 = T236;
  assign T236 = T2[6'h27:1'h0];
  assign T2 = T3;
  assign T3 = T237;
  assign T237 = T4[6'h28:1'h0];
  assign T4 = T5;
  assign T5 = T238;
  assign T238 = {T252, T6};
  assign T6 = T7;
  assign T7 = T8[7'h48:6'h20];
  assign T8 = T239;
  assign T239 = T9[7'h48:1'h0];
  assign T9 = $signed(T11) * $signed(T10);
  assign T10 = io_signalIn_imag;
  assign T11 = T12;
  assign T12 = {T96, T13};
  assign T13 = T14;
  assign T14 = T84 ? stored_Weight_i_1 : stored_Weight_i_0;
  assign T240 = reset ? 34'h100000000 : T15;
  assign T15 = T81 ? T16 : stored_Weight_i_0;
  assign T16 = T241;
  assign T241 = T17[6'h21:1'h0];
  assign T17 = T18;
  assign T18 = T242;
  assign T242 = T19[6'h2e:1'h0];
  assign T19 = T20;
  assign T20 = T243;
  assign T243 = {T246, T21};
  assign T21 = T22;
  assign T22 = T23[7'h4e:6'h20];
  assign T23 = T244;
  assign T244 = T24[7'h4e:1'h0];
  assign T24 = T25;
  assign T25 = T26;
  assign T26 = T27;
  assign T27 = T65 + T28;
  assign T28 = {T62, T29};
  assign T29 = T30;
  assign T30 = T245;
  assign T245 = T31[7'h4e:1'h0];
  assign T31 = $signed(T38) * $signed(T32);
  assign T32 = T33;
  assign T33 = {T35, T34};
  assign T34 = io_signalIn_imag;
  assign T35 = T36;
  assign T36 = T37;
  assign T37 = io_signalIn_imag[6'h27];
  assign T38 = T39;
  assign T39 = T40;
  assign T40 = T41;
  assign T41 = T42;
  assign T42 = T43;
  assign T43 = T50 - T44;
  assign T44 = T45;
  assign T45 = {T47, T46};
  assign T46 = io_signalOut_imag;
  assign T47 = T48;
  assign T48 = T49;
  assign T49 = io_signalOut_imag[6'h27];
  assign T50 = T51;
  assign T51 = {T60, T52};
  assign T52 = T53;
  assign T53 = {T55, T54};
  assign T54 = 34'h100000000;
  assign T55 = {T57, T56};
  assign T56 = {T57, T57};
  assign T57 = {T58, T58};
  assign T58 = T59;
  assign T59 = 1'h0;
  assign T60 = T61;
  assign T61 = 1'h0;
  assign T62 = T63;
  assign T63 = T64;
  assign T64 = T30[7'h4e];
  assign T65 = {T78, T66};
  assign T66 = T67;
  assign T67 = {T70, T68};
  assign T68 = T69;
  assign T69 = {T14, 32'h0};
  assign T70 = {T75, T71};
  assign T71 = {T73, T72};
  assign T72 = {T73, T73};
  assign T73 = {T74, T74};
  assign T74 = {T75, T75};
  assign T75 = T76;
  assign T76 = T77;
  assign T77 = T14[6'h21];
  assign T78 = T79;
  assign T79 = T80;
  assign T80 = T14[6'h21];
  assign T246 = T247 ? 18'h3ffff : 18'h0;
  assign T247 = T21[6'h2e];
  assign T81 = T121 & T82;
  assign T82 = T83[1'h0];
  assign T83 = 1'h1 << T84;
  assign T248 = reset ? 34'h100000000 : T93;
  assign T93 = T94 ? T16 : stored_Weight_i_1;
  assign T94 = T121 & T95;
  assign T95 = T83[1'h1];
  assign T84 = T249;
  assign T249 = PTCount[1'h0];
  assign T250 = reset ? 32'h0 : T85;
  assign T85 = T121 ? T92 : T86;
  assign T86 = T87 ? 32'h0 : PTCount;
  assign T87 = T88 ^ 1'h1;
  assign T88 = sigCount != 32'h4;
  assign T251 = reset ? 32'h0 : T89;
  assign T89 = T87 ? 32'h0 : T90;
  assign T90 = T88 ? T91 : sigCount;
  assign T91 = sigCount + 32'h1;
  assign T92 = PTCount + 32'h1;
  assign T96 = {T98, T97};
  assign T97 = {T98, T98};
  assign T98 = {T99, T99};
  assign T99 = T100;
  assign T100 = T101;
  assign T101 = T14[6'h21];
  assign T252 = T253 ? 24'hffffff : 24'h0;
  assign T253 = T6[6'h28];
  assign T102 = T254;
  assign T254 = T103[6'h27:1'h0];
  assign T103 = T104;
  assign T104 = T255;
  assign T255 = T105[6'h28:1'h0];
  assign T105 = T106;
  assign T106 = T256;
  assign T256 = {T258, T107};
  assign T107 = T108;
  assign T108 = T109[7'h48:6'h20];
  assign T109 = T257;
  assign T257 = T110[7'h48:1'h0];
  assign T110 = $signed(T112) * $signed(T111);
  assign T111 = io_signalIn_imag;
  assign T112 = T113;
  assign T113 = {T115, T114};
  assign T114 = T14;
  assign T115 = {T117, T116};
  assign T116 = {T117, T117};
  assign T117 = {T118, T118};
  assign T118 = T119;
  assign T119 = T120;
  assign T120 = T14[6'h21];
  assign T258 = T259 ? 24'hffffff : 24'h0;
  assign T259 = T107[6'h28];
  assign T121 = T122 == 2'h1;
  assign T122 = sigCount % 2'h2;
  assign io_signalOut_real = T123;
  assign T123 = T121 ? T217 : T124;
  assign T124 = T260;
  assign T260 = T125[6'h27:1'h0];
  assign T125 = T126;
  assign T126 = T261;
  assign T261 = T127[6'h28:1'h0];
  assign T127 = T128;
  assign T128 = T262;
  assign T262 = {T274, T129};
  assign T129 = T130;
  assign T130 = T131[7'h48:6'h20];
  assign T131 = T263;
  assign T263 = T132[7'h48:1'h0];
  assign T132 = $signed(T134) * $signed(T133);
  assign T133 = io_signalIn_real;
  assign T134 = T135;
  assign T135 = {T211, T136};
  assign T136 = T137;
  assign T137 = T207 ? stored_Weight_r_1 : stored_Weight_r_0;
  assign T264 = reset ? 34'h100000000 : T138;
  assign T138 = T204 ? T139 : stored_Weight_r_0;
  assign T139 = T265;
  assign T265 = T140[6'h21:1'h0];
  assign T140 = T141;
  assign T141 = T266;
  assign T266 = T142[6'h2e:1'h0];
  assign T142 = T143;
  assign T143 = T267;
  assign T267 = {T270, T144};
  assign T144 = T145;
  assign T145 = T146[7'h4e:6'h20];
  assign T146 = T268;
  assign T268 = T147[7'h4e:1'h0];
  assign T147 = T148;
  assign T148 = T149;
  assign T149 = T150;
  assign T150 = T188 + T151;
  assign T151 = {T185, T152};
  assign T152 = T153;
  assign T153 = T269;
  assign T269 = T154[7'h4e:1'h0];
  assign T154 = $signed(T161) * $signed(T155);
  assign T155 = T156;
  assign T156 = {T158, T157};
  assign T157 = io_signalIn_real;
  assign T158 = T159;
  assign T159 = T160;
  assign T160 = io_signalIn_real[6'h27];
  assign T161 = T162;
  assign T162 = T163;
  assign T163 = T164;
  assign T164 = T165;
  assign T165 = T166;
  assign T166 = T173 - T167;
  assign T167 = T168;
  assign T168 = {T170, T169};
  assign T169 = io_signalOut_real;
  assign T170 = T171;
  assign T171 = T172;
  assign T172 = io_signalOut_real[6'h27];
  assign T173 = T174;
  assign T174 = {T183, T175};
  assign T175 = T176;
  assign T176 = {T178, T177};
  assign T177 = 34'h100000000;
  assign T178 = {T180, T179};
  assign T179 = {T180, T180};
  assign T180 = {T181, T181};
  assign T181 = T182;
  assign T182 = 1'h0;
  assign T183 = T184;
  assign T184 = 1'h0;
  assign T185 = T186;
  assign T186 = T187;
  assign T187 = T153[7'h4e];
  assign T188 = {T201, T189};
  assign T189 = T190;
  assign T190 = {T193, T191};
  assign T191 = T192;
  assign T192 = {T137, 32'h0};
  assign T193 = {T198, T194};
  assign T194 = {T196, T195};
  assign T195 = {T196, T196};
  assign T196 = {T197, T197};
  assign T197 = {T198, T198};
  assign T198 = T199;
  assign T199 = T200;
  assign T200 = T137[6'h21];
  assign T201 = T202;
  assign T202 = T203;
  assign T203 = T137[6'h21];
  assign T270 = T271 ? 18'h3ffff : 18'h0;
  assign T271 = T144[6'h2e];
  assign T204 = T121 & T205;
  assign T205 = T206[1'h0];
  assign T206 = 1'h1 << T207;
  assign T272 = reset ? 34'h100000000 : T208;
  assign T208 = T209 ? T139 : stored_Weight_r_1;
  assign T209 = T121 & T210;
  assign T210 = T206[1'h1];
  assign T207 = T273;
  assign T273 = PTCount[1'h0];
  assign T211 = {T213, T212};
  assign T212 = {T213, T213};
  assign T213 = {T214, T214};
  assign T214 = T215;
  assign T215 = T216;
  assign T216 = T137[6'h21];
  assign T274 = T275 ? 24'hffffff : 24'h0;
  assign T275 = T129[6'h28];
  assign T217 = T276;
  assign T276 = T218[6'h27:1'h0];
  assign T218 = T219;
  assign T219 = T277;
  assign T277 = T220[6'h28:1'h0];
  assign T220 = T221;
  assign T221 = T278;
  assign T278 = {T280, T222};
  assign T222 = T223;
  assign T223 = T224[7'h48:6'h20];
  assign T224 = T279;
  assign T279 = T225[7'h48:1'h0];
  assign T225 = $signed(T227) * $signed(T226);
  assign T226 = io_signalIn_real;
  assign T227 = T228;
  assign T228 = {T230, T229};
  assign T229 = T137;
  assign T230 = {T232, T231};
  assign T231 = {T232, T232};
  assign T232 = {T233, T233};
  assign T233 = T234;
  assign T234 = T235;
  assign T235 = T137[6'h21];
  assign T280 = T281 ? 24'hffffff : 24'h0;
  assign T281 = T222[6'h28];

  always @(posedge clk) begin
    if(reset) begin
      stored_Weight_i_0 <= 34'h100000000;
    end else if(T81) begin
      stored_Weight_i_0 <= T16;
    end
    if(reset) begin
      stored_Weight_i_1 <= 34'h100000000;
    end else if(T94) begin
      stored_Weight_i_1 <= T16;
    end
    if(reset) begin
      PTCount <= 32'h0;
    end else if(T121) begin
      PTCount <= T92;
    end else if(T87) begin
      PTCount <= 32'h0;
    end
    if(reset) begin
      sigCount <= 32'h0;
    end else if(T87) begin
      sigCount <= 32'h0;
    end else if(T88) begin
      sigCount <= T91;
    end
    if(reset) begin
      stored_Weight_r_0 <= 34'h100000000;
    end else if(T204) begin
      stored_Weight_r_0 <= T139;
    end
    if(reset) begin
      stored_Weight_r_1 <= 34'h100000000;
    end else if(T209) begin
      stored_Weight_r_1 <= T139;
    end
  end
endmodule

