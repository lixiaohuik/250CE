module AGC(input clk, input reset,
    output[18:0] io_G,
    input [18:0] io_Vout,
    input [18:0] io_Vref,
    input [18:0] io_delta
);

  wire[18:0] T107;
  wire[19:0] T0;
  wire[19:0] T1;
  wire[19:0] Inside_G;
  wire[19:0] T2;
  wire[19:0] T3;
  wire[19:0] T4;
  wire[18:0] T5;
  wire[18:0] T6;
  wire[18:0] T7;
  wire[18:0] T8;
  wire[18:0] T9;
  wire[17:0] T10;
  wire[15:0] T11;
  wire[7:0] T12;
  wire[3:0] T13;
  wire[1:0] T14;
  wire T15;
  wire T16;
  wire T17;
  wire[18:0] T18;
  wire[18:0] T19;
  wire[18:0] T20;
  reg [18:0] reg_G;
  wire[18:0] T108;
  wire[18:0] T21;
  wire[18:0] T109;
  wire[19:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire[19:0] T26;
  wire[19:0] T27;
  wire[19:0] T28;
  wire[19:0] T29;
  wire[19:0] T30;
  wire[15:0] T31;
  wire[7:0] T32;
  wire[3:0] T33;
  wire[1:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire[19:0] T40;
  wire[19:0] T41;
  wire[19:0] T42;
  wire[19:0] T43;
  wire[19:0] T44;
  wire[19:0] T45;
  wire[19:0] T46;
  wire[19:0] T47;
  wire[15:0] T48;
  wire[7:0] T49;
  wire[3:0] T50;
  wire[1:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire[18:0] T55;
  wire[18:0] T56;
  wire[18:0] T57;
  wire[18:0] T58;
  wire[19:0] T59;
  wire[19:0] T60;
  wire[19:0] T61;
  wire[19:0] T62;
  wire[19:0] T63;
  wire[19:0] T64;
  wire[19:0] T65;
  wire[18:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire[19:0] T70;
  wire[18:0] T71;
  wire T72;
  wire T73;
  wire T74;
  wire[19:0] T75;
  wire[19:0] T76;
  wire[19:0] T77;
  wire[19:0] T78;
  wire[19:0] T79;
  wire[15:0] T80;
  wire[7:0] T81;
  wire[3:0] T82;
  wire[1:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire[19:0] T89;
  wire[19:0] T90;
  wire[19:0] T91;
  wire[19:0] T92;
  wire[19:0] T93;
  wire[19:0] T94;
  wire[19:0] T95;
  wire[19:0] T96;
  wire[18:0] T97;
  wire T98;
  wire T99;
  wire T100;
  wire[19:0] T101;
  wire[19:0] T102;
  wire[18:0] T103;
  wire T104;
  wire T105;
  wire T106;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    reg_G = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_G = T107;
  assign T107 = T0[5'h12:1'h0];
  assign T0 = T1;
  assign T1 = Inside_G;
  assign Inside_G = T2;
  assign T2 = T26 | T3;
  assign T3 = T4;
  assign T4 = {T23, T5};
  assign T5 = T6;
  assign T6 = T7;
  assign T7 = T8;
  assign T8 = T20 & T9;
  assign T9 = {T15, T10};
  assign T10 = {T14, T11};
  assign T11 = {T12, T12};
  assign T12 = {T13, T13};
  assign T13 = {T14, T14};
  assign T14 = {T15, T15};
  assign T15 = T16;
  assign T16 = T17;
  assign T17 = T19 == T18;
  assign T18 = io_Vout;
  assign T19 = io_Vref;
  assign T20 = reg_G;
  assign T108 = reset ? 19'h4000 : T21;
  assign T21 = T109;
  assign T109 = T22[5'h12:1'h0];
  assign T22 = Inside_G;
  assign T23 = T24;
  assign T24 = T25;
  assign T25 = T6[5'h12];
  assign T26 = T27;
  assign T27 = T28;
  assign T28 = T29;
  assign T29 = T40 & T30;
  assign T30 = {T33, T31};
  assign T31 = {T32, T32};
  assign T32 = {T33, T33};
  assign T33 = {T34, T34};
  assign T34 = {T35, T35};
  assign T35 = T36;
  assign T36 = T37;
  assign T37 = T38;
  assign T38 = ~ T39;
  assign T39 = T16;
  assign T40 = T41;
  assign T41 = T42;
  assign T42 = T75 | T43;
  assign T43 = T44;
  assign T44 = T45;
  assign T45 = T46;
  assign T46 = T59 & T47;
  assign T47 = {T50, T48};
  assign T48 = {T49, T49};
  assign T49 = {T50, T50};
  assign T50 = {T51, T51};
  assign T51 = {T52, T52};
  assign T52 = T53;
  assign T53 = T54;
  assign T54 = $signed(T57) < $signed(T55);
  assign T55 = T56;
  assign T56 = io_Vref;
  assign T57 = T58;
  assign T58 = io_Vout;
  assign T59 = T60;
  assign T60 = T61;
  assign T61 = T62;
  assign T62 = T63;
  assign T63 = T64;
  assign T64 = T70 + T65;
  assign T65 = {T67, T66};
  assign T66 = io_delta;
  assign T67 = T68;
  assign T68 = T69;
  assign T69 = io_delta[5'h12];
  assign T70 = {T72, T71};
  assign T71 = reg_G;
  assign T72 = T73;
  assign T73 = T74;
  assign T74 = reg_G[5'h12];
  assign T75 = T76;
  assign T76 = T77;
  assign T77 = T78;
  assign T78 = T89 & T79;
  assign T79 = {T82, T80};
  assign T80 = {T81, T81};
  assign T81 = {T82, T82};
  assign T82 = {T83, T83};
  assign T83 = {T84, T84};
  assign T84 = T85;
  assign T85 = T86;
  assign T86 = T87;
  assign T87 = ~ T88;
  assign T88 = T53;
  assign T89 = T90;
  assign T90 = T91;
  assign T91 = T92;
  assign T92 = T93;
  assign T93 = T94;
  assign T94 = T101 - T95;
  assign T95 = T96;
  assign T96 = {T98, T97};
  assign T97 = io_delta;
  assign T98 = T99;
  assign T99 = T100;
  assign T100 = io_delta[5'h12];
  assign T101 = T102;
  assign T102 = {T104, T103};
  assign T103 = reg_G;
  assign T104 = T105;
  assign T105 = T106;
  assign T106 = reg_G[5'h12];

  always @(posedge clk) begin
    if(reset) begin
      reg_G <= 19'h4000;
    end else begin
      reg_G <= T21;
    end
  end
endmodule

